��c      ]�(C ���e�Y]��@�5EW�}���e�����6�C ���(A����WX�5V��k�s�!�]8�Sq�C ���3��}NjjT6�bc�)��'*?�E�_��ՔC ��F��Nt�Ի�Jsw��K�+��C�8��C (���.�u~$�u�Tb��{q�R�JA��y��\&�C Ʉtl���'X�T��V>�������g|y�W��C 
����~�v�Ҧ�2�	�\��3W��89Jvz�C `>h�ρ7笢�<�BR���i����٤�[ȓC S�2%ԽAj�R���؃z{"M�i�B�\�)vD֔C �:1�f�����c� &�ht�]�����-��dk��e.