��c      ]�(C O�̐����ף��ߧ����u��[rM�}�]�C ����B^�V�e�:��bw�t}&Y�ܶ�v�C ��4*��ô�!��w���l\w+d����d��{�C �4�,�/@ ��������;��9�q�4
+8�-�C +i�W0�8�W�����1��pu�#ٿϼ<ĔC �l7��o/ؽ����bs4Nqe���x�הC <�����KCu�3�C�ɓuJ����B����C �8�S?�C�f����,[o��<����S��C �*��������Bh��31'��[Ө��S���C t�"֮��MKt><Sf�>���$�zc8[ףq�e.