��c      ]�(C %IZz��z�=�Q󣿑�B�����+y���/q�C 6:lT�!�69��f�zU��b�Д.��cŔb�C �����SY��A��U�ך#�|�{-�d!�Gug�C ��~[��xp��ǨJ�Ƙ1��}���x�(�ϔC "��$]�1�#hͥ?c��d�!�� �E~T0�C ��1aG��A���Y$�a�����|�<�8e�C �N8HJH�ҭ�z�����l���V�<g�I���C O�\�O�yc	/Q�֘I�bCh��_Q�.�ՔC {P*h{*e5
f�h��k��[����%���_�C �ʳ��bW�P>'C(�Nx/>�SU`���e.